Library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

Entity FSM_top is
Port(
	
);
End FSM_top;

Architecture Behavioral of FSM_top is
	
Begin

	

End Behavioral;

